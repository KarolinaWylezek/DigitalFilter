LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.ALL;

ENTITY REG IS
PORT(	DATA_IN : in std_logic_vector(7 downto 0);
	ADDRESS : in std_logic_vector(9 downto 0);
	CS : in std_logic;
	CLK :  in std_logic;
	WR : in std_logic;
	RD : in std_logic;
	DATA_OUT : out std_logic_vector(7 downto 0)
	);
END REG;

Architecture behaviour of REG is

subtype int is integer range 0 to 1023;
signal addrs : int;


type storage is array (1024 downto 0) of std_logic_vector(7 downto 0);
signal box : storage;

begin
addrs <= to_integer(unsigned(ADDRESS));

process(CLK, WR , CS , addrs, DATA_IN)
	begin
	if ((rising_edge(clk))and(wr='1')and(CS='1')) then 
		box(addrs)<=DATA_IN;
	end if;
end process;


process(clk, CS, rd, addrs , box )
	begin
	if((rising_edge(clk))and(rd='1')and(CS='1')) then
		DATA_OUT<=box(addrs);
	else DATA_OUT<="00000000";
	end if;
end process;

end behaviour;
